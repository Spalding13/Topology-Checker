******************************************************
*auCdl Netlist:
*
*Library Name: HBM_testcases
*Top Cell Name: test_1
*View Name. schematic
*Netlisted on: Jan 22 14:09:27 2015
******************************************************

.INCLUDE /dummy_organization/projects/users/amit/testing_thesis_subcircuit.cdl
*.EQUATION
*.SCALE MICRON
*.MEGA
.PARAM wireopt=1111111

*.GLOBAL sub!

*.PIN sub!

******************************************************
*Library Name: HBM_testcases
*Cell Name: parallel_reduce
*View Name: schematic
******************************************************

.SUBCKT parallel_reduce GND PAD VDD
*.PININFO GND:I PAD:I VDD:I
XD1 GND PAD net18 sub! esddiode areapd=2.925e-11 perimpd=150.00000u nf=1
XD22 GND PAD net18 sub! esddiode areapd=2.925e-11 perimpd=150.00000u nf=1
XD7 PAD VDD net1 sub! esdvertpnp areapd=5.85e-11 perimpd=300.0000u nf=2
XD17 GND PAD net18 sub! esddiode areapd=2.925e-11 perimpd=150.00000u nf=1
XD18 PAD GND net18 sub! esddiode areapd=2.925e-11 perimpd=150.00000u nf=1
.ENDS